module Memory(Clock, address, Resetn, data);
	input Clock;
	input Resetn;
	input [4:0]address;
	
	output reg [15:0] data;

	reg [15:0] Mem [31:0];
	
	initial
	begin
		Mem[0] = 16'b0000000001000000;//MVI R0, #2	
		Mem[1] = 16'b0000000000000010;//#2
		Mem[2] = 16'b0000000001001000;//MVI R1, #3
		Mem[3] = 16'b0000000000000011;//#3
		Mem[4] = 16'b0000000010001000;//ADD R1,R0
		Mem[5] = 16'b0000000001010000;//MVI R2, #6
		Mem[6] = 16'b0000000000000110;//#6
		Mem[7] = 16'b0000000011010001;//SUB R2,R1
		Mem[8] = 16'b0000000000011010;//MV R3, R2
		Mem[9] = 16'b0000000010000011;//ADD R0,R3
		Mem[10] = 16'b0000000100001000;//OR R1,R0
		Mem[11] = 16'b0000000011001000;//SUB R1,R0
		Mem[12] = 16'b0000000010001011;//ADD R1,R3
		Mem[13] = 16'b0000000110001011;//SLL R1,R3
		Mem[14] = 16'b0000000111001011;//SRL R1,R3
		Mem[15] = 16'b0000000001000000;//MVI R0, #0
		Mem[16] = 16'b0000000000000000;//#0
		Mem[17] = 16'b0000000101000001;//SLT R0,R1
		Mem[18] = 16'b0000000101001001;//SLT R1,R1
		Mem[19] = 16'b0000000010000011;//ADD R0,R3
		Mem[20] = 16'b0000000010001010;//ADD R1,R2
		Mem[21] = 16'b0000000000000000;
		Mem[22] = 16'b0000000000000000;
		Mem[23] = 16'b0000000000000000;
		Mem[24] = 16'b0000000000000000;
		Mem[25] = 16'b0000000000000000;
		Mem[26] = 16'b0000000000000000;
		Mem[27] = 16'b0000000000000000;
		Mem[28] = 16'b0000000000000000;
		Mem[29] = 16'b0000000000000000;
		Mem[30] = 16'b0000000000000000;
		Mem[31] = 16'b0000000000000000;
	end
	
	
	always@(Clock or address)
	begin		
		data = Mem[address];
	end
	
endmodule